/*module Instructionmemory (

input [7:0] A,
output reg [31:0]);

reg[31:0] memoria[0:255];

initial begin */

