module adder4(
input [7:0] A,
output [7:0] B

);

	assign B=A+3'h4;
	

endmodule

	
